library verilog;
use verilog.vl_types.all;
entity beep_vlg_vec_tst is
end beep_vlg_vec_tst;
