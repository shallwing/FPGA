library verilog;
use verilog.vl_types.all;
entity flip_flop_vlg_vec_tst is
end flip_flop_vlg_vec_tst;
