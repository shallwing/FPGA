library verilog;
use verilog.vl_types.all;
entity saler_vlg_vec_tst is
end saler_vlg_vec_tst;
