library verilog;
use verilog.vl_types.all;
entity decoder3_8_vlg_vec_tst is
end decoder3_8_vlg_vec_tst;
