library verilog;
use verilog.vl_types.all;
entity encoder3_8_vlg_vec_tst is
end encoder3_8_vlg_vec_tst;
